/*
   CS/ECE 552 Spring '22
  
   Filename        : control.v
   Description     : This is the module for the overall control unit of the decode stage of the processor.
*/
`default_nettype none
module control (/* TODO: Add appropriate inputs/outputs for your decode stage here*/);

   // TODO: Your code here
   
   
endmodule
`default_nettype wire

